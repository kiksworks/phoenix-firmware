//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 23.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
iunkIMZIuocjzH7zkWmaZEpngGJPqviXSWcUzerXqX8iun5LMoYmS+phMc1wZpq6Y99H4mY0f0C3
j0uw2dR8IZmatv+2AFBiSpnBxuIofPLKthmPteQk+5+pm6gow4/5b6ivErNs34VdJ5CDaQ10oHcb
krzqrTXsh/u5p5lyYyDu1Burk/kz4ea4c3JgIC4of2UOsb80ixnmUBvCn0M69XXt9MRk5DWOvdod
KswF/QY8eCYFN1Yo9E2Rc0HPSbYYqlcAHNLsIX4vVGA5fW3ZbLgaH7In0Kv87ne/42LIdrXMtwJn
ZTGZenwC3fN8HRnzzmoXGDg4ZY7jGgw7z6t38g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12704)
TTABDGrtnyA9oQRJ9buvZ66JmUi5dzk3ah7Ou1ukBc+klY578ppw5ztFKKBZ1bDv+AWSeuY8cGMV
ht5HVQ3Tqpr/swLGpbXk6OnvQUCC+K9J5SM2FqxINm3iq+Vjow10sqzV5x6yySmIK1lZ+IMeBAEk
iH4+3+NyKkSvW2QSfpE5UL1xC3heHBYvH/Rr09zbJKDeHRsPRxc2hNaM3W82STZ7BUREs/Du/JMM
+MA4scRsqdhJE8zzQkVKrnyp2HhKRUAat68NnzFRkxqBthHtQs9n3tVj8Bst78bYtdFrDWh5cA3B
/Xwpkv0L0atUheEbTOyfRubb9ABp1CoYXCI/HILZ6iTJKtvpkMiIlBKXD2mGOekWyx8WPfYZQOuh
/cgvtj5aqoQAGO8McQNkIGju/mDZk75qHpcFtl/4hu+YU7AVd6IrnbwkCtypwetoFQhvip1NDxs8
dnV6iCZGr4DNZMsdX7cWIw363KXijJnqpkBph0Rui/zPJwEgXPPvx2C1VNgsZyUcnAWz40xYJosI
JcU9ymYYXbOTcs292cgZIqnzkaqFOqsoW2qxeUHUnDiNDSyYwhf99CX/N/3NG9Kav5ryASx+4Za7
wNRyIOUuglNxQEvd/EJJd5NtXNzIt8tLKE3pgG36SNXiCnNvkPK8pIwmEj7ZLlW+bAQu3iCNtI7E
8GP2NMPbOrYjXig3owE65fsGywwSrCd6tH+K7oIN7+KWCf86NLZznZ8iiXfXiqM4ytXad7BOAi5h
A1JjL8pQFI/oO5L23WlFlDl7OoygptJ7wo7gTTW2Wh8NeG0VFn3c22JELPLds5f1F8HxYpf9syPr
xIT463I8I2aW9zKPOKwqJ8kTDEs6uLAx88xFY65ft9NkN+m3w9sBMBMRNrkuepZ2kh90p5adMWL7
JO8DMtTQXDNVUncW7Wt6IkTiC4yjrXKvxAAsM3wltHRWQXdqfge8X8NTGsJ7iHZQlIjH32TGdd1L
sndWB75s0gRM0GPQGWe1JiLkMbDIjJ//BOnciQW/XHTqnDr+i35IadT2/LYg6OVBe/SagQ06h4c5
56XXLvKu4vZoPqvu99oV/qn4zVSistrDH7EuSuVRPcyeTvZuTOWovcBuS16H2UVaKMn1J58YlG6g
RussQteHUBTJ+UEFGi/q1tJY7HvSo1Y1hlChuFr94oJg/zU6P7PhqvjrhYn4KreSHTcyKKJdHS+q
iz1WVkP0+ck9Nvj/phTsPJnkZld6f0gnZ9CVzq8uhYpZbQes5f7DjgeSQCcYBlY1x9dccbufh3ZT
+rR0nOnnwjL2Uf3h/EFWDYgFd5KxqDU5kmm4h8M6EifkGLwNOGDUxC+Ngc1crT0/tKtaXRc28R4B
SzpJg/MhX9WjgAgEqSEJjSZm/PQemPtuXTPsSvcstXvzIwkVDvWCuybattPGsVn4juPJDTlaX6O2
mC2wd54qkcsIj6sYz8hGxBOnji8v2WxfVOPwgzHeHCAA4LKL3HwxQMvUEroWa1NwaijDAGx6l99Y
KSd0o3GjA0cOXqStjAF6Zn5EsNHKHmTo/N761Twq+zxXAfuaPqx8wwMH+02pfU0TmP1puflfaBX8
/IO2HwK75Q70wlIjjrF6h0wq19X8AC6nxylAbMrA6BlX4gJ3Gidd7c3I5LQJ9ktJH4xR3pGyoUpJ
/HqWlB6B+bko+nqqrOa/LGO4fltCcT8VEE/+N4y1iyESzKbQuWAc/fGexMxaX1BmcHHuAYymQzzq
OHHR/5EknDOOoSLVjX4AXvW1D998O3LQPbt65kA3uxHeaHfeY+LUB2w+F87QIGNnkiKdWSdF6Fuf
1m0xyRaBHEsq9se03aNEqiU3cwIvIeYpkqNFhZM1A7ckYhCXdZ8g/tC2nU6S0WaURHOpkyf9i0li
mUOc0NzHbSxgl6sCwp6GcS/CRWDZ+k8DRxKjQFu1Un4kJw6AOn9ytd1JMqT0+o0iSg6ZvnFox89m
gRv7hYW02N2mnt/qJHMrejWZHndI2yJAxb385D853plFlpRFtTAczGsT71ciO+6taun3xQHLNu4R
6I+c5F4J0xKSJ0U8R1szgwLg+FtG5SMNBqJP3QuNzNhKY6NS7hg+m1BDqckSsEaMNFsmwnnKHy5k
bRYjcPFCSY7btFOOOI8mbkU7HyJxiI3QtOWwEGwY/+cOPMVOpB7W7dNM5IpT4149FUZiWnL8g7zq
atKabvExbbTiLVlWqepZDlskIZJxErECWcT+fSmGTeWXcx51KPPLtHOJRnPVjw5gsKXLt4mYRnxK
ssJ8bZgwhqWUZs9dm21zaev6yI7MOBeFCaPHtiOVixfGsqVFZDUvxngoKbOCXWlpKqi5OIwVIcmX
4okTE1m1Krp53z6PuLJO95Y1WYqcC0i/MR05kO3Bm1xzW6lKwES++smKyitQlFGIjvxwKPSI+SrA
zR4ReN0eOMTgutupmSS2WUivqckBmS3ow7iCFRpxz13YqlBvJBYs5wnSEHgqjqs01TN7IgI/FTOZ
6RyWjoDr9zv/L4/1+7SSyV2FBiqwxJk0EGUcpD1fZhYhgROanc0KJImNz+W8uXd04mp4wvcgz2Or
uM091FzELCD3Nc2ZbPUJAKgz9KUH1Msb81PfNtxGeX6zw4l60niOnR2tahewf1WxeV6RY7nF/mL/
wZC3gn5bqGYrA31EhnQu1pilyOv2ge3kDWTOy4KZdZF2SPRQfkAZln87x/hTVM40zrcrORlO9NC1
KoH5vmf+FQq3qyF4pBAoLE64/kGQGSsNgVeIsdCslbI/HyfkPaWCa17WIIQjJdD39zp77aFPudjU
/w8mTk1dH04YD8UcPW2mEBgqgJR0wCgIcL0YP9WJJDevVogvhWSOMNkeJaVbOb2/URLN8ZhVqTWP
JUP9OISAiR+RNZqB+gQGTWze8YJS/MnYN8I3DgmCm9+Yex6fFWWVQ2Tccb8LDB7y0zXY3bCYevSh
h2i0QfJJjL+u0rU2F3+wQgiVw5cwo+5MySEFdXy4pb0zlT6NMAO3Tv3jH+nkZegjguVUWU7bhqB2
c1FuUG6rtoEpNiY4ldahDgC45gLkr8ZyPxtjpgzWBpkMaTs7vGruZrgoDPRrIk6caomuVlsqRk2w
N1KrEEFx6o3ZD1EikMLxysOJJs+X+6ycZigVXhzERLmj2bAgzeJTfNs1CCKAe9ZPGWJSC7ckG4z5
I2elu0mQGR9ktU76g38YRrv3amrlHMjNzLFsMOkGR2dmrLmowS5QjHJzhZ7W1d8K3+984BbQ3U0G
QgJYgPRflmR9SCZykNDdti02lPpAvCAny7qM80JOhtL4ze/+MAKHBCnjKTLku9ImQGkdyMBuvuUy
AU3nL1suBRZVi/sUSDp8gXHpHG/OR72p+sYdLRLcAvRPqHCt1le+smpWJIAHtMCg+54NLgUXaUsc
VGfFYS2alX9X+M3wRjPCiHhO6GJ8GO8NOhpbe234dbefOd7OylyI+NJRzMTkepvuIKt9zoK4khMS
sfkO8GOCVVUCBdrSToD99Pq0OPhKwINEogNfc/bzpvNKbGGvjtGhepyJV3Tmw72+DUZfnaqEmC8x
6yIDDs/jvhJGGlUhJFoeJ8/qv2ZgsZ4xJXUr9JvcevFnUqNKiQnFy2cwuvkbhplmzifczmwfr08q
GPyW6DqQ6DD8HGnLsq3vGPrAiLER43wd7mzUD0ZhoVJZ4Z6C3Ppy7PsyEFXDnzDb1aGhLalqUy2p
alAdpCuMDHPqdHw62tsZmRAyIb8f40AkI3iNZltCqkxhWEh39+SoHVAjlJGlnmayBq0xZrq5VsxT
zhFTjAsCLHC1jInZQmnqVu5TfKqa9EG2O6H37amewlp75wKyOjfxrF66cEtI023tmKLLneIjKSYT
8ynWIAZmTGOH52BfXPdKauCJi/UqnE3/VQq1eQMWfqbDAY/zxAV0QIsVNpP59BO3G213BSMwdNfP
gYZPy8HToJCiA2jxeJM3wyBj4yE7E4OI9SS9wAUV4+LUFFcwr7+nStbQxDUenm6Gg/k8u5eHCvx7
Ggm+7+jgM8mFrZEqYVTms9BoIP6gT+52orupGDWk29Tqz8oRDDyHA2tVd/xaNy1OdLrCvHzikNI+
8reA/nY9WWFZdVhb2n7a1Z7Dvu1nB2zuCJNp3jU0k3rnNme3pjIcORE76iPs7/cN2pFAWQXQc4Nx
daZ4t3gmBKc2QhbL8MTr0FtqFS2E4hF88iueNj//8LA+u3hsYEgDiNwdqau89cb69J1uwbHWz4KF
95i4gMdj56HVl7bdm5SRscUxxiCFXu5KPGI3iJSlk/6HrLxg/uuqLJNlDXVNXGtImZygp4iAPP70
/TQ9lRTpOTi1DHDPwJC0HaOerQREcaUr2jj5bOOrqknj9XT1BAkWEOrzWQUUpEu1y9v9wCxhm+9i
Bjs3g8d7t1hQ2qcEeoag4lTyeeABP3JydB2uhXOGtKtqdeDn7gjO6931tXT7VJInPQRJwNgCP+Gs
H2iUUaSgl5L/eZqMPXGT+Hq4tRX+kZWqQFNpH7rBjvl+3mj4nfveqjulycwx5o7AGtUr/EZmz74C
ndn5GfSBf75UcKZYtwFUQ67XlgjkZ9PWqeULt6JCE2LerOiz41qHKcq0fXH63EO+h1hsbiaKxSzO
l+Ej2jdUlgUZXnHpnOf4HzPUBg3JVoKTtHcJOHEh8hLKamLsQ8WvCs+4exBdj92ET1net7uK1pgX
h2BNGdOfvuTjDCVUflFd5cYXbFUcxHma7c+PzdZstMq8mK6wqucebNj9Rm06/MDLK9q+Puk+NuqG
9s5ZjufoETRXULOyMuqeiC4VW0rDEDwwD4C9Sl6ttXNm2BLR7OfKFpSXJbgQr7ZltcpzKDsNwqW9
zKTHorqQ/mxLTSc2cwsPqsJlK5ZnsmuswukUguUtcMqGXqkY6MkkaeIqFhO/Yyy8bjqBexUmhpBw
vKoxxpPV7zxt0uj6vRchhFHZj0RDajiMyFTFStiyMjqTEc9iXVh7Mq0hBgJa2JkL8eM4387ERg9p
jRnRKD2biEcT+DwuZxKItFcgyIyqPkELLkzXr6m4k5kIk7QlfAWKX9VLE+k+AuvBFubtsZ4go5Ce
kQll06VY8v6IKkhOs/AyQvEQ0634LThXtkKBiYF27ATp+kMK2LyyVUg7b9Y8m+z4FEBjiFut4G6p
fUpsdZ58t8efYYiobkVRnPEufIXfm1KjSTeiV2E9TAA+3O0BHyfz5edjgDQru8vYUXhr6PdJEXH+
HeGdA5iXwr3ZVBUmJdS7FiKkQfhy+u9WefXxh1lccgELBVx246JPHLV+UbWLurtAg++iTqecU2KP
qMnBA2nE6H4XrlXKjcwwxWolL0BBcfWA8gi8NEIhBo4yp57fRaZMkk7D+VHTvjhnWP4SL8R/wg03
39cxrrcB2Rb4vy13+e8bolqjqypMfQEcG1sbObDP0TjJmYtSEN45tFEayzp4171MqRidUBJ1m329
OMyIox01z8f7xOanbiaOfNAkWU8zUqCV8XdsYDytbYdbsEjC7Wvd2O3jTldE7BV3b/26YpuRZLco
kyjmEASDyEsc8FnPNxFlpeMsEezvsQkzhNeAgd2FHi+SXjsJ4S1c1K+xCugdxMiL8IwWgRK+W4dC
Y1We9kyst3I03vLRXYy5/JYjxWScHFrFlus93chuTglSlib5NPlz+xJDNwBLYfDw/uiTY4h6votC
uHHFO7dj+xOvPEXjlqxD3fBibxM/800WzyaILU7KUSGFKlkLJIPhEW/wJ+zyAUsoTlAqwUoAqdeB
OHJepv7zMV1I484YWHM+eKuLL1BrHmNul7FPI5QUAbPmbKqLAHG2GDtZ/GUYbtCxCSxLnv9nWgFm
Zq4HTpjRcYQj2wHrX/i1AxzA0fcdZatTwwguDrA23oBBkuTl/45Np+2ser5StimUoQa9d/qZzOr3
oMLCF3JPDqBqawQLisgRVEI65QFwqDsL4R9lCpMiE/M79jxTNUaNs4/DwroNHtqAfeXvYhC0AB9O
FIuUXbhttzVIVEYJYZoxmnSYS/CnmYfLctLQoNoCNxTi5BDjZ+UfgXCmqZOKWdN8/8FtjWOfT/PV
sxcea5WAnf4JyvPn0PEV0GB2v15cd7Bxz+Z35YgKh1MLNjL//syKufTDR6HaOHAoobTu/HV4ppr/
1F/of9GrjRfbnbTDZZd+HDs93INKLU5mxQlQ40z5zxJrQENN22KtRfbU/Y+ItCLS+cTw27qngvLU
OPBYcZyrBuGFVPK30P8+74EbI1LA8z/xn0ff/tzA8iCU7gU5bfI9C5kGL2baZABbL+fvYB/2v6F2
AQt8ogRctWa/0FYev2e0JzqrmTrRDgcof583yqk3uiywhPyihC3+c2cyk2FJUqXX7vIWLNHaTMrf
LrZmV2bzdw9v+z2u4LYSvk+d4g0BXCh2gxUsLmIaLSUcFGs2v+20lO9L8qNgttITbAMWC1U9X8w1
o3HkFg+xmV/78dY/pn4EGXVV0L+Gm7oR/7QbSChuwKLcoT6/w0cAsAx7LjnOPqxuuQD/X3wIPnjR
YRxCLZNjaujOoHcD7UNAuDY6IsfHXba80a7v4gb7dlH1iOVKStZqJpQBnq6g0h5MD+ctnGgdpi6Y
X8ohawRECeqHRyizsHlCIg74ey4Fu0hkkZaw9yH6bv6FpshER14SpP9WX5XZ7LDsSUyilhJJQEtv
nUQOFPPME0gcWwMD3h4zFvDrBHDtrIwS8Dp83TgDJK/r9e0onokZ/z16bDvtm5KeKEaY9BYW8Z4g
mU/y6Ia0kEe5HC2kn4fOI7LgQNfdCMa3U45r+TbVbYa5GjPumfFxt+2qgsauUFf0xURYIhYNZfDU
GHeAz5fTdLUdkoyypEvqggrT7dVXSF26sTMXuPkgW3eyGeJ6vpVUPIv3MLX4En6guIXwB1rxKTW0
5kr1oA3tEbCz5dR7skfTe4+eiI/sow2r/CEYs0K1Xu6quvJv06SPHhW7LnjenBQl+TsFIJD/v8py
kMgGyVLLaCPa50PWRsRol7B3yN8Hl2WmMFL7HCrTTZIJcg0hWdALZBQlotgef3NLvWhCBIuecgUO
3fWNg9yQxaKvwsvIXfVtj48vqjgO6yeIeawmhpwF1fwIFFJlqRWqacnB0E1/gzUpbHaBfkoJNApl
5qrRBTPElmLAJeMobDsXq+AuAtxyDvS/AAG0+gTerHTzmG0Gobu/eK1KKsqASeA7VzuaMi+9Luwd
c5niZPOx7XVY4r13FY2TYcYUrwiuCj0TS93zwcxEHZxkkJPCDaxCQqc1l8PgXr1Cqd7Qu76hMZsM
HD6xMX3f3a2NZBy8yg2hoo7Iqx9b7UW1dmV2gKnwi0KyULh+uvgoMmnXov/C0FzpJ11rcBShadXV
NBMRbSOZ9KoYW55SCMbcM7H8Rnov7Dssz4aJi4O3pOgkWNQlI2quzncNEnmQTeUhJ0RZ/uaSkYZs
k3IpQsNQBn1LQPfde9EgIkKBjogvKopPIt9FcONNWG8hWAiUtRF+wnZonmyHt1feCTVMMYi/bD/M
oNCctxJCU+iemxh1jMDBV0JTiLJ/EB89v+TvGPuN5t+QgRHsnpNmDooUggC7hyWPGHNycUqsjHs9
MnyF6m/v6G/PGHRwtubqnYmlFHWhJKbCOtZrENBBKoIK3f39nkzp/w3N9i6c81W97iK+XjbAD8Ge
hYVtWvRFcqQsmZXfcc5/3dIkpvj/ts4uh7vSIulZ2ZZc12xUN6H+TqDYs94ON1OkOg480HiX8cGc
DpinA8AWt2Zi3QIjsdeGDOifTKI1SSSeCb3+3Ej900XMHN+21BSbwMOUMxt9t20hY2pAtqw2omx3
iEo3uBlGnL60XAbU3N/ucxVdF80y9lAyeh71zHe6/+UrlbL5nZqgqULM21plJUeqOACNcSXLY+kX
sEIy9P1/qTFU3oMBuTftMeeHC8UjK2XkateHsFqpiYG4CTs6SbhIYmy938Qdi2ayHSiVaVHyBvj2
+fB954m71deqp5E5h0TCa7J0trsZ5KGCg3eI6TrWTCohYeUmMpQ7W9oes9gdC2nGP+U0Btic+sF+
jo1UYCgGKnm2F3hb9WDdLFfjmKpjjzjGRYgEuBa6DpaX+HxhVdszlUnjOHqoPqF9Fvqy1WqrB5rm
RTJmCbT79MFgh4prpyPWxGBOqQ8StlFrzl6oNrIvRqacaA6azwyNkoPTeOiROt3oUrAhKqT0UvOf
MHfZ1l6sioHHAr4+tyspvAY5IM9giiel7EudrUUK5aKx6pw51IGxbhIO02yyOJp88rjmV8X9oa0E
tZ+SQQ6TDHmp7a4UdimYAoHDdkF+w8hs/CiTfMJC6IHNrFpae5EhhBmWxdMDXYA3i3dtl7A/WoMQ
1P+fmYt32T6wJi7/Ewq2XAAU/sKH8ZL+WFcdh8QLHTsHfrRD2Pap6OrGXuAOtn7BQ4wixxrFw4um
hNqsfGgYt3FWauAYbOwgZyL/YhReMEd4kT35SoA4UOvqj4N+ITvs7JgqmBrX1FKy9srRQFffOD46
kcbzidrYlvwJ1vDY7FMqGJDas6MSwAak/XdbU+yytg8hkOtpr8xzbxAiJVGjA5uA0ulWCtSsSeNV
krH5deeCaZ5MXaskDGxFwFS6sdsG93nq2FGKTm+yCzAlQ/VKHQ4FL9AXF1NFLHM0f2SeXaCmkX+E
ij9wqCWY1nMnAOPqhD71I8hRYhNLoyrLb47+vtYg7b7Efa3XXeEq6uUVNGyfRfZomTq1C1D4AQ1a
3irQD7PDZ/BMYiKWYVMgb34bczww8wtDRl7zbHoO2rg9akFaFh5BdD4WYTcUqZkVIG+puU9gCQ+M
6hdRuX5Lw3DIhJfZAVUvvjI9ajHKsJnSyEU4eroocNbQRosyd/Mb0eta0TPhVMfeysJ30CEh8X8h
wbMsnAz/k2pXXEhBu9sSBK5NyK3u3FK6DcWQ+WKISU/fYLLcGDIecMUKo2/Pz3kpxGyX+zeyvqNj
26fmKxRa60w9IAPTRowoj9Qm/Q7x41lLqw969Mp0U5lVPagS+5UHKRc6ZRggoSRu/m593G1T5Aq5
/EaOv2xBrYaYVqKZfWHozNQbbCmRPUtyQOR04a1lLI2dnK2uwqrmJCErvmLqWn1Ej7wUznPvukDP
mO0b9+6sk3QGJ3kXtWAXQtTtfdApt9aQuqSemY8DI/JTvSzawvH2M7P8F8w0wu0WfPMXUxMlm7Gr
WyNnTysyPI6QAkGY4o3PLsu1e+JQpFDSJ5X/tmiI0yo9qFO1gF4msqRnzA1ZSXfq/mM+DwLr5WQ9
4V6FHu6mykGjSaLKgUxHl51EXZDZ9SXL2+DmuGfyjOx5gtp1J1Tec5ikMmPdS/2IlmPcLDMk199c
7KhlryDAm1REP4xh1V7+JU/ZowGgmiWHh1vX3VxdROUi4/o4G2USXvwZYk8KFBTP8yKb9AIyYXb6
C3awfRL2lbHul6NFqLoOonPI0TK4AefQXbhvr0ag7EefBWFn+Gw+UuUOTnH9KDxDIxx7c53PITiZ
a9iTjX6Y5wiWB5xq94sWDRPtzh/nLlN2hGTxeBNRtRJ6muLjkQ+g4rinsODgHgjhaatuYcrwAp/1
rlrOwkd+XdruLaVd0loSOGgnUWlQ8tBjgfQb4fQhtWn/TXLtCScZVdElttRi/sZS042ZjGscAuW6
m2XSABlDz3M6ylIL6q80Kn4yr33vscQYnu5n2VJaddOtSYIYwy81eMdmJ4Wqq1D2wfK1pgn5q1bk
nIpv6qjR05c2cqkD+9qRfrNiJRvthEn/rbg/sKrfeY453cAsN9ZUVxS0iJ7tvWBKqilq3FYwmAOV
zVBO719azXDAxXdGHKJdSYOOz/zBN8TipxDoFWHtDeSk0nSlUu3WkFqL2xgg1awCS0m9YJeIpJWg
jwyM38/eLtU6PPza1OjxcI6aZKKZeqwKcViJH0nzwMpRdSEJB9rfjtXysfeudc9/y6b/vV17Br+Z
jK4S1anikFf0EzRvOWuAkvNDxmdsF/ZEnunjqf7LzGn1uUq9CLM8mgYCBZT7Z2f47VmH0JeiDclq
XrTnHvg5JJME0+gaAE7qOe8O1dzzIsIKr3LkzR0xoawiLp47SLmYUUwtVoN0TXAL0RAoNfexY3Cx
slBDKNf4MHYe6h7fekNqLoL8ElGjQqxy7rOca8p8dn6tPQ7o8crxoG1FcKHB0crc46jeKkwIQA+L
Dz4d4zaJbGh5WAZ1BmYFyyGsyA3Z3TF7nggoI7mYPOoOfPJWTIJgV4TetadHHFFza6rlmhbWkOsn
rJNZ4k89Phc9KcbhYfsYrs8j52oJ5e2UvNCTYKt3LLmRjssiImdiDOnrDhyJ/MTQ7sl0zgA+5lrC
qfpBuMP6+cQVgmORDZUqGI9viLpJ4aoaPyXgYYjA5OIMkoMK9bRWC5ppcHFcjUk9ZJUVNMYPknhU
jAv9tXOMzenakcITkGS1uGfzCVqtuFv2IglPgX7eUQ2P4nFo45/JFDPWprNMiQNdFyFQ6V5d3iah
EYvsNgokHVvCrOUmnMKcLOArqq4jWXB/zW9tL62ISQI/a/P6jgYJZuj83ONseqW7q6//lCg+c30q
B0vmXwEXB5M2KK6tsBb9QPMMP0F1kPp6hfR8hmgdNZMJYaDvPglFSV5iVcrrSV2o59KuUILD9Nur
psPAoMS9lVR9h4Ct0a7etfrHOkua5CqJS0XzgfoA4sVOHGfiUTTLb6p2xCM4DQI6JmrkngB29VJy
b3AX4aihKAwo5ENOfqW+ZeDGNZnX8FdizIuMHSG3HVQdr6MmY9QC1yzpRZnSpF0nxPlC/YATpqvA
I7LaFvv9xtMfPwFD4MfvtbsiU9WTB6xDjoLHvUdo07McZ2Oybiv0IjrnbAvsn/IRajiOHXxvej3O
8UfwgQ3f5KoRim1cLe4rWnBlF5d+Mst0UvePtMBJFa1DeNmC5odTp3x2N9bSyHAJPpX97Ork5Ewp
uOQYhMFNFYHZOAyuaXqxwciokYmeOYhUFsEC87bTrvUCqCCEUxEh5+a0ycbbgGzJWjl3eXC1fG0t
DbeZTFd4qpuv9CXaCTRxBUGhMtN8DJpde5nSebErpsCjg4TZaoaJ0551j2+brljSj2Vmzo9bMOVX
8VWLjpvuACALwcmlFwfUqgzqXDwDkeh8JcP1A+Jhcx8Q2bEsG33OMq7gn8i+/IEKTIsdTjxb4ng1
MGKSkdF1Yt7VmnYLKQUKLaPdnzGrHwo/hJdluIlvyKH32+98N8MmiqezJrdozqBLSWw1GA4Alq3h
N//TYpMVCH6QMwroH4RNEQ86oU91jlcrrb08OxsLjHW+qdfT9grw/NeRYckYsaAID2EGK4PoE6mO
ttHrAg3X0qz5I2zjNYQtMaXVdkxZ2+LP2txvp1Ia0i8FEQp7tXdx1LmFvlLtnZ5KzsgExMm4BkXi
gmD9ZY76FUbs/lfbEGqkNM7wkGdn61MhA6IknIh55fs3APVCwEG2z/kTb/0HFTVJYEzxD23136Py
5rZS9nzAtyEjncpFnhIiELyYFPUz5zckt0tBdILH+8BovwSJSMLytEMt4YDs7tTxsTg6zEypv6TU
+Ha9HW7UlV/4fX+t+RP9qWkLGGSCm44SsRSbflTzXDu7H43yvRC7rNPxQR4ocHwRfpOziToJSFn5
qlNUjPjwwPt+CnPWFWdn9b39PB7+vw/5KArXXSW6hgflex9EFRjBYDJANT5t109mEbwHXLb0z9tV
bNnfzXYbZYTmd5efWFK8ABi1H/J8/IzW8WIZLGgSHLIgLhB2MOFazYFOoLvvAvKR4P9N62jtAQHo
TlaDkx3PJx7wadFo+cdUaglNGCYYmB1UaGQME0mNvH9tQBHJBnhFsTkaZKBDgZKAqe5dQ2fEgsZX
NEkbH2kzzYZSMFZj/jlvElDZvRTa4FtXQCo1J9v8remQGGBriDb5KjwshEaPB9SdbpBIkcDumlmg
shh5eQK5S+TMgJqYSl3j0rIyPKSc6xwhcXVw9I+BOqFt/Ko8l7O/N302dZJhmKTvo/xGv0Ugb3TD
7wUoT51UQubHFTlaW65edt/aY1BVfcS5+M2LQeyLk8ITgCwhNDlxZ/13gfHsx6gTxl+iQotd/KRP
4+ydI2q/c8TgYbEROsyOI6t9M+N+yEB3byZninnf77ljI9wwZjI8pYZpwgIByeEaaMTpyXkGk/W/
7uZuZ/9U30SeojQG328HQ2DOnGPEMkxeY4NzIkBnIfjdwd+v9KvCmaorVKmw6DXnLYl97oI+JDJ2
uKmvoiHQvmvSTzPL4S9evwEV01so3W1MAiMQkmBeK2ngVYoik38Zv5VyyzIejmHTATJOmDlmd/hK
if1O1uhV84nDm6YccrwR5D4XN4fcEi+P2KUfecrg8frYoVH40uNkvJYS/5ANrTZpGkT34JqRUgE/
TTfYVR8deElgml3YcMdY/qyRXRLoBnQ5ruyDiqfRUB4YilIsBJSNU8uryyc+ZHiM5SJ3FTePc56O
VIpqYaB2h43zrZd2e5Gfn+revj3jsLOKqIt7XqTV7OvlkoiP9XsiJ7e6iy1nHbLN46LwDA0M4fkN
QJeyEOHTYQ3wKE6S5wzSXnaepOr7689dlzZ/zlShO3Mf5siDXqwZrcsGWa07GzjEQ6hDm96VJxil
+YNLRIVEOkNtUalWG7Ew+Yaq1C1eEv+PlGS/JU7MSv+gzoU3OqdpHEw8SIFA6TNxopvSXNVZCLy/
iCv1NVIg6lGuAY9MK8LWusXZAoQ/geC5YYfVHDW8AfFGUHz+rMMEfQooy3Bt78kmWxUt9QtbbJSi
NvXa9B8vaZwdRoktJ5GeL7cFXV+NC+/wtJiJd9tkc98HgfoRX4JSRlKmWiXzVulQhNb6i15aH5wV
5VdE3JJVLxn21CK2KdzhsSadVHfADjgMaJE4XTYDjz+7YPCO9xvWDm8wiwWBSRppYBWMFzIOsjVU
MItxa8z5YT46PQwI7LEqVmyaUBokHhjlLkGlQGq720uorlhcLMBzOqy0HyznkBDVGig55iOCoLhD
slbQxijmDbZpyJn5ciTO3U8CQpOtp78Pwdlqa2s9aom1kL+7t0m8X/ipQcac3aC+E7RaRHPuAMFV
hhox3csX9fQnGSk0pw9AGAiiLMFzqzSC5ZnCC0ieQNmlYN34nccSSj7SIp7x/23Xfw/o8xfSsp4O
eskNfxye9GV1+riee1O30jpXUUGXZJGe6TrdKBT/6gKg21XAXYw1sJb1O4thDWAqrz6bLc8m629D
B174mCcMNNmFv/EcLIXEwiXQnPE3rRhEfVy2XTHM8w3cfBaPj4GT6WCg6k7fxBr7i33yXFnAILKJ
57qDIhrs4T86EYvOFxjBHXbplKyChZIJb2ZR/sIn760wbeMsgeuIExKNduQT1bLhZg6OofDyt0ln
Vvt1QyC5sI8RxH3t9vHq/Ey+0R3G3KMeLhQOaib+DMFd5InaNwcRMONvXTHsCGHyvEjBCFD65RVY
uMT8wR0khC0XWEJ6QJEB4hmvasN6i3t2f/XI1nE41IK1tEJ5b7cbbnlkXgKa6D18RR5nXRs3dgQx
Yn485fDWki6bXIFke/pnaOcGtHBpfGdzapXwKzCU3+Y96WoFIGmBgH+LLULhyLpAT/zTYEOwDj1c
EM5aBbCujDBG8ETrScIlG6v8MBLbh9Pie7L7OlHKZMSWlHbO9RLhtTI6ukZ9Y2txyVFMyuQ8izgT
tXjjhrOoWh6FnOeJgmYp1xb5iCbMlx4uS7/9ZOZjMHspMgr3zOXatTNXvAxUVPWq5NMUiS9RdASa
+VwxcK/ns/zQEzoIVtmeWbcPU8d63uZp2ZuDYIk5EkHLfqZeVlJGCghksG8kAfE17HeIVHes5Qj8
vLFaNXJq+IZxzgYZXnk0xR8mRp0LmBC2Z7ewIAZ2kjGTwF317ntO0Jtoor7OVNPpMKRufVzdTQIl
ASmeiCQeWma25xchKjg7lhK/VMXMzdMkv5/kIrCxlTlBLqWbq5XOao80GADGjvJfgVfyD9LzCLjm
o2rAfghMBh0v4edeYs2C/u32PXaO4mxTb8IptEdjbVzThCoB+69MuSuYFa876MKUbY2OjVK6p5Ei
c6j37/QufaKnrWHgPT4fnBtEMovrkHCvG7r+DXle3c8UDZzFGKIEllDqGFJYmDtYzOtZKY5lhfX2
7uRoXbrKoHi9IR1/wBp+p+OZnDnuJmF2qnPLbDxy0wyTKwCjuqaGd3+T71JPUFw5fZrXa1nz1Y7Y
+anbupn3djidn3GWXOJ5atKmrvbmXBdUD+UAkTYxXOmsw5ZwYUV5b5D5HnJrOP3+1ZChuHwVriDk
MwMwnvRshOn3USnZQG3bqJlsPRG3ce9Nmr1kzFL7TPT86VP1exMvpN/056jt8A2uRM9+GxXE2+Tj
fXEF1UTtEfAFJ9FetPxbWGwuFcfFax2OnZuzfEK+WPnZ0VIhxz/BC9nH4DxUWcUtxwiIOypHybS9
6+1vE5VkyAcbgjSMg0YHxNifwAW2cssXPIpGxwTwl9tWZomgGLTqdEmGYdMPaOSU2ngblAsfIRbO
/jroVPMEne1ryDptICBTG1fUxspxwRzYRja4KdYG4AriWZSHSUqN2fcdwBDgljC2MfI189Nnhi10
EcJMV8Oz7//dvuLhKmNaKdLh8oXlP8+sVeGCuEsf4kkwsxUuRjglVaO7kBzw1T79RmyiyauiDjVW
W9s/fn5ca8x2jJfmpuosGO/4ddAqZ5j+s9ku9ovprMvF2Uey516Z7J6VZJJEqfBKHzZhVUsSPGE5
mcGiyqiQc1Xab5rIUSc6Pb0A12daV0EUeoj2pPhXRRNE1aCxeKZ9oPQUo+ql3DwAaMgMLg+grzmt
fgreZQ7w/IL0dgGaYdg6hWE0Jg0+5Fr4SHX0bvp22DjCrOtO6BNZvxtWL0fbC+4bZg1rvir8T1sD
MOSgtANrxBcp61x1o53Nk7nAst4CLo9nelUuuCEThWLAZk0aLk1hiAILBqkhMF2i/cbikplQO6hF
TdIdEkSRZROMjsnsmMI0wfs4ZAggROmhkbhHIs6fx64EXQeQMzOG8GCN1jE6mjcQOfCiwHe70BHJ
LSkPEQq9eteQj5PYGyrxGD+Sa0oUPnIqbSMA6Jj6dyEkjzxaDGwusgjMDuqxiBpG890RXVdjU8IK
74oWrWQW3fOjARZ0k3YFky5G+oBsTjhDDXWF7I8fI1CwBQPIMO9gcIcbVtlWFHZngRtQPBJQohMZ
mEYGQnKra4txdrRHD8PJRvmbS6f0qsiGEdYYnNxZYtCRzPO1Jj2TmH8Hog4iIfnL/ZG16cMetldv
eQLfY6lrSzOQZn0CooM68SLKneiZHTh4EcWgQxaT5BT+ZAX7XI03VsHlpvtiGFJIBszNuVFI2CwN
UaDGZA7HmmijeTXRudAmlv4l0dXjq0UZBsli1MRs1Ih/lc9xS7d9NhKaIX2WJ0Nwfq+r9K5rUH+7
yoYUWN6YYd2BBiyVnwzSVYrOV2jtMoilB5LyzppK6l9j/pMEV8cgWhAll3kfhXbiw+TGyr1kPHve
oNW6+vsOW7pO4xcZ+WpJCA9F1tKj7EX0O5J4iubL8MnZecJVnRalhOhcnGYRt4NkcB7uFI9Kbzjf
LgcfUFzQYwSzghkUxA4DA2PSFGtphwa9HyAY61xCHwT6hX4/do8X6RE9SJAKvxrGCnOQjoPGfbl0
YHE85BOIuqDuDv500lb2jfUQCbxDwTn+n5a+8z0BEvsKCTKTjQgLiyI1cs/H2kyV4SRNolLouBra
pGl9+4RkFI8SB/29e8JxzGFWx7ympWC2pTx+z3ANuIpeOj5o8VYtPwkEbD9PO2Y1UV95+v46iHwY
g8nKh8OZPSIMH34aKwfvvmCHRyH9AFqfGjIzjxsapiUMJl7hTMb9nx0ULpVT7otJ/6HpHhv0irTD
Co23FncQemTAIStfQjUQcUWCplVI2x+XcfbbU/O0yoLa3Wun/3soolZW/0ZMJlh4VDhqFbLaZ466
IdRAyoRH/5YqZ72AIqS1bwVP0i46JSl3Z6wbu6OzKriIMPPnlTyCI6MZ0LZ8WrbF12UHNxaP4ZMb
aqLvbQ0TRiUkf6YatgQ3jMFwgbcdfPws0hdGl7/k1CfqrXxB7QhUm9IYcN5r4tvwe4rSXp8SOFHr
DMEozcFbyPBWDeoGiEsT1Oe5I0EMS4N9r2t9S6UKTpg8BaShEHd16MO5+zqDt6dK55pXjs8UR7KJ
ExnaUMNLNEJ0egFt2p9Omm2PsK6POpKcrkCvvEki6MNju5uezo5Lseo9SqFsgGoYGNJ67QIPMPB+
Ntds0nXd7ZyyVUYlc4rST6+ZxVU0MOSfwBrRXm7I70YA7xHZFe/bUMySJj//52xACzeGWhfoVCWQ
mhVxpghbXFt8ugW1cMe5v18p8SzF56WCZ1bORl8ZR+IWTJDNfyXQNOPwxQgOGFDhYce6xG7a5+mn
EIlHWIcg8aRsYOOAwh47AGEqG1tpDATGUZ4cHqDeI0744tjYl2RpuBJWNo6fI3Fn1pZYqKkNmjqr
985zEhSpDhzqYi3D+hYAhmoueJidXuMYJ5V6sP8RIiVsfUfxqgZw1wY+F8fAnV3YJsdJZvvll5qI
NpHETjZ5YT7t4odnaOPRpNqt9psHy8usMeZ4XglOgq+NztcUx57c4HH/bWZDxNHyUzFFUxe8nt70
jpjP3cFhjY6OoYiN91xZdPblISbt35atGP2iAm0EiobBMzziltjZguyAqAppv/6s0la9VXCXI9IL
ft5ZBT6o1o8FW9ihG2eOce3CDRuV6cBGSywYslgKodFZmuUsxJLpk5B5aMeAokoCKPlfmv1P0tm+
sUe7gyM4KIXgfzUeR3Dvxj2yM7AKP8e/P5+ByunG/RF2gZdlDviKw6dsct37oZLm3PJaOZlQcfu/
pRCZhZ9G+V/NpdJclK20jlZS+FkJsSSilkJBxG5yAYWhHn7/bxhbvrZESGJ+b2IKGj0=
`pragma protect end_protected
