`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hT6rbQ3rOAUV8nMPbrM3W0IRHAdk+2E6HbvR+eo7fIgR9BakZolH5K7C6w4j7zKg
cdN4njEBe4TsALX/d2bw7T/SGMTmOX3m2LRG/DSKbKk86xUEc6m219fA6TW5VrPs
s3KAasYBTaEdA+g+eU3OusEN3y8nH+Z7AMvWj5bC724=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12784)
K87fbEDQQpOqNfnwxNLPVG/rQS/VSjr2GoB5GFHF3FfPVmQTktA6yp+yzKwQ5abN
ANXI436Nkh5BslChmDSIAzyrpKDBxyDTxM/FNReUfDmtOWpp+1vHa9+pz0nFU7k2
xLBA7b2WwU2ylaa6503geMIUWJgn1ihmDlGwMbiUrnA2kBpejI5CYBLRF/cpITmO
aseVuqnmpQ4XrL8t+RhCfRbiZWVgiHagET2USDcP8lpLrdN8lrtniqDUsj2zPJNw
38h9gzZ5E8Z6wqah4/a5FPMKl/NV5UvBs3nm2MR5547iwc0PfYjRrkFsQ8OyDE6U
+WPciNgTKoLskSf0+M3t8ZrQU/QNKJKBUb6wPs6r/EIhVAwcC9uAib5Sj8oMlXGs
QVKv+vd7UFzkyYONtOz+JxgkT8WLZh5Gr5y2PAMRk2a5XFh8tm4V1huU+Lcm4gk7
DNs65T1k/STb61PkFAO6pLvoz80hbUIYMdFni62ik9DLGlHQG/nTjZwITLKftRii
YWdbm6lesbDovdTPrAKryjI5LHicBxGmu/PsDj14Di7qfjVAuUDQrIhVx/xtg20B
b86i0NRXWEkQne63O9VUprmoHJJu5Z+nL8VsCeNNQc1/xvd82rCqHGi83neSyCdU
EIsgxMqkzvMjut07fvPQnwSJuqcdqqAlX3BAIfIvC8OUUJUcOU9PNrHMI34r9oZj
5IYPiYZ9CIQ6ScDfUuD5zU7qMu3flmHliU7Zj2t4H0yC81IY+1IV2WD+Nvhzbmai
mcP5fVQgC/Aa+c4Ij8L4OkJSMqaQJs7relyprg7ojlNLF2pySSbWCB0gE/ldkFAe
RAhaQOF8uiDG4Tv9Kl/46JehBqOEwxW8fF0zf6DhUp8EVcIw3UdnNzAMLMrwzOsG
zEOo6LVIFXbsHr/Md0mOBlFUtG9u113q/yBRgUwf7s4PwPSTWyXVar8kc9QfAL3s
oKMH+EYd+ev/IuTR7btmSHwSEWFlGudMwBo22URjFDtccWA7n3hze1kaCGOgJBED
tOXn3s6z9Es7vaIuDMvuGG78EIOhPVy9LDtjbgq/GqU3xqbDNjYsRRebCxBm+OII
kdELuOaC1I0Sgo411abdHNrTj33QkAXclbsuKt+JrszxL4DCJY1+tzn27ZOQmwPR
7OC87ag6kDpDcHqyhF581amHdszvyok5Bn/0zNtqzvASJQct73zZYFKsd+xP41Rs
XcZji0IAXI2tFb8gEga4ELbwioQ8bTEjMtKQbhu7kni+uIOu8S4eXAzZaAJ0xo5n
69im1Lr1CawXp2vL9JmuYSUwG+1p4vPXe/oRmy+DS6j1pTR+dDF4rFjJz/REcI9X
Y/kqjV7OdDemXp5UDz0SJFkmfOcIL1rG8iAOc+k1BwONBkkJW5IR7m1ilirlFccO
H3osVkjGRqruAf1Bk5TlQ1cNrg/cQro8HI3jba+jPwQzGNmMB0deaAumd2V07e3Q
qE107y2lj+TUh4SHrVF+E/M5VJxewTHf0eGmniXeMWMwENfO/Mnk0KjpkGzP21Ua
fth1fZgpxngBJTJk/zAsUudy1BcBPOT2cN8Yfkbz5Hboid89VsMTasHzgs1NcbnM
wIwZJRClZ3ngaUafidEh2RVV37rJ5ZU/c8Bqfu0GUCJy1oTyQVXgZ4d9XdrAJVAT
naGU4QrEzFWS5I9PA8k+ofv0wlutucC5gWK9F8HHXYl8gwcXfNTABojvStWteEZP
7sdtYv7NufgIMy8qT0433JQyCRek0dvsngGLEfkQ5R3XVa6Ve25EamMAC1qfwaY4
PiL2WAAPmbu/OjNT37jA8L9HM4WHsWw2WZtkNfO+X1wElaFRm627JSnromSY4L+B
RxEZkXge3BE7TDvsQsRsS6cAf85dxilTQG1h6AWwN0aoik2qoo5Qt1TS1OUfOobl
6isqXN2BN2CePQoNCmvUeosQSnGJPvd271s6c2/zhhv4CgGyAc0hRp/kfGhxnh8M
SiIV7FS2HchWUNtKHALZXi40huX4P83UQyglLCzRX7HOZIIv0yNHTtyDIVK14sIm
9csq3/4gpI9U9UDGZOnk1QkU9Oixghizm5Y+tvE822zTTur7qK5EGnyRjU+LI1Gs
fAgIPQOg2xj/YuX1fiPJ7g5nqNxseDQEXOVARyjrJOkHKh6t4W7GhfSWNPA+ZCip
Gqf+RkewTB9XsYdSPajmOeH9HkX/sKnrSRS2cLQNQyNc9195Q2KtqXRCBYltnUdk
ApIp9dwAG3WSZLNA4jMkCeJVrcHq/eubdpcWHGUAnFMyrSY/CNN/X7+bMQz0cMmD
45V9bOdBLa1nWlyhkXpuoky2/3JOKbW5ls4RVLgcg+Rw/tsrtNZJWM1aAIEtNliG
BxOAOtdgsDf07qR/bP7KnXhikVzBUwjRfGp9/cKpofA2SAziekM6ythMz1a2ogys
ydh/rkDcLAZa101g7J6qn0jw6ugCKxN+77/IhTY9owmatxRowclCsASzKk8Et14l
6sW9kvJ3rE+lJ0tiRkWxU0rCKQ99iCcdIL9hV0NuMK2La5s854wKnwfYBT39l6Fg
+RnKkwrsL3brZn5m8ZXAFR4GS+65pshRMQ86Jj07l3mBcGPOBPEAMlcnVFDhKwgm
/VeHVW5L7DUq95XKi8PjY9oKER5bG/4GYov4UZ3PHdUuAmzzeJWC8y/Vwie2Dcrg
ZcmxTzT+wKukQTwD5cPe8kcmWX6knxHmwmFwXDhTEOTIK5bYZuoBDEXg2P3wA7GS
jqVs/LeCmrOHptrIDONisVERKcOJFOSX3Fz4Vy0AXH9U/drtWfn3JKXskzsyvquc
FCca3CeHsA4Kg2pj0p1EkKKa4KdnD9Y8q9F0AHCEiY6aVAFdtJcoo1jHdI2NNKVU
yJtIxB1ybphvwmfPu5zzuSR5py4Cj9l/77bOUp5bKbcvWyrmHsJbAC+Hs+FE6xua
vdbYQEZXKOw5bSWtaFbs2MBD6Wxeho9fwvovR5i8rf4uYtdl8LmceJR3yiCod7Wc
0vNEYX+9wmRiQxau09kepC/zUfxslQeuxGIgKD7NPhVMOIDu0B83izXalbTwLvXd
FzayBlmVJgk5jV4BCJDq/+6zhkbZZ06wQYfg7PlWpzPGZcBpDAFepq4MzOhpw9LF
Jtk8Z2kI96RxFZis/kTcuWndXy3rmCF3JmnoCKHy7cmfhyuTVeEI4JYXF2shcYHD
DD8trh35r4mQjscFGDk7aF97kaWiJ7v+dF/3RvG4UjcIGkpFsKKCGhCgR9elYKe8
D/pK722NbClgBs2dIluclEXU4IYiGJJy6mtdQa4jeNWhzOMYF2+Qj0ug5WI51bDe
Z1fzB2G/4ge7uGiiuseGXFhAMRVZj07nsmyR3XtFTaNGj8icaLf9sKw2A0KwiLtj
GqtAOAgcdRb/6jBYUUilk61vhUhjGknbPMHq1Cv6RS9h0Pt0PvWOdQshSfBBZbEC
vzz45YormVcCMXuKrBihnaxmX2kdnRFQbSqQANxEEUOC8bSfgD1jmeR5JQ/9ydpi
EaP3D16njSy4Odvmmckd93xN0PEOFCeTnCd3NimYiQU9FdlYrQ0e0RSGgWq+rS5h
Iwt4nCab3zfAPNQvFNJoPOepVta7I9zU1H1lOqQyQKGHQ5079exsVATLO8t9U/+R
A8fijS4GUZwiJoULC3uGtfowCVQkMdLC9X0r6EnYpwpW5HdfCCT9sWFqh0NSd76D
vrkb2B5CopRL2wMsk285SnVq1XMY/6kaI5E6xHeC/7oZQhp5dXOtPQXgy3hzsj7x
M243CExpbdPrdWPDH4C8C78grGRSDfoUqeXodymBHl5Sc9BKFIRB4c9IgKSOcPEI
IG3hLcRmmesIyuDt7PEZkpfS/y67J3JIusDyziihMGpgtdFtirOFgmESYS+B6sYi
uZ4bK1dEIf5x+tCzopd6XDz13DeXg/ajptHPtVU5ZpC+cTbLRDOG4p4X/ER0oFOl
GU8W8OiK9QuXQ65CaMboAK9BGq7+t2PsVCHlOAbWnz19sVcvn6mQZyWvmPvI7Rrk
1REv0sHCtYiWfcKLXm0YCWFW/KPPs6Y85vaR6jmUTXfXH9YK21t3fPtX1f+K1zVR
lrlYJpUe6V5/LxD3rxW4T5M92JlxlReYO4odTY5whDTWT65N21HJIkzDiuBD965/
cTgQmu3KGhWi41covDpqfHNJZJzJqmyl7nTl/WaMg4mAJLpqGrCpBpd8LUlQgoP3
1ag34WYTLosvmgT/srGEbFnJGdQ9cWBmCm9dCKtouTo2oBe1EjZ10pCiVAbC8ULW
z3xI+7nF7/SDZgSDXcCyTl2eWAoPUCGWggga68wnq/b+9Bnw3syrHUsPZ0WYysgg
Xu/oCU6/I3Xkdeay/IyRrouodTf1yHgU5EmLxhg/LSCuvoGSk2C0J30Zlo5cS+8F
sedjEv0DEi59bLbGMeEafZlkW0ZUIxqcR8fO/j3HQEp+DSudmRlyWhx/DukWHTAI
4iXQqzFb4nz/5XUtrF6W9GkkqRkuCZFVCCtVYktuqmtWA6wUe+Dyaekkvwn/ow5D
z/gHBgkLaLVFclFdp4E1PkPIbGPsgU7Ol5Azx1DaOZKtUOfZG2xh8+b800uV2UGA
OzwmHxwmsUfKoZgddc1dudChXnGbd9AoausexQ3UyuR9Nz2zqTPKKoDUCYLFCU7Y
9y5H4GHKPhjFH4027rVtsaQ7c00qevCxJzjtp1MXxjMbWVDPpbDawVd4GXtB/xr7
NM8noP+Jsu6JZtQAHW0cwz725TMpqXAq14dy3Ilz+X7wqs3T3Iea2NHyQIRraVD1
bwDIAPn5dWIvZ0lPS9YhiFVAP5RjxqMuXKGFN826/eNT4cj3QNHCgNAPE+NlJuny
M9VwdUUxdYdngXPaKX9DwQZLC7uxiJPql8vvsLGLvc1/vIaqej2rKEQdv8DcV0FA
95gF6F+v/5Ap7QAq6sRoDWVQSFCGZsy2nkad7PGKRjevYdAmYU8G1RYkuj6Qv9j9
UCoJmJhP7657UJAUUiWgIxZbSLjBu07G60v0cKuu2AJrS4Bphd+Gp9EL/JuGS0nv
N+T9DfM4x2ghb5T9rbPmSIb32CecDKXm9QI8G2UmVdKpHLeKQ9U6T8sCXBGYq+Tw
/S8/9sPdcV+utd4mEwgI7pQRhuIOUtZRgq4flVDDl62XXt/dmSO6wTERQ1tHXwhY
JXTI4f3uypWiCZUIGGrJ2tK4kG/sZO/VOGfGI/Xn0KJW7uM9Brw4Cz6Ln3BT08sH
cMwpmlUnpMFSyyC0/LqG7QsX07Yh0/+WuB6l34X616UFYPlG8DztD/WLXw5o9cpQ
yQrHO65HDNTgGttycGZ14cgFdIK2avRfliDJ8BlUkMXW6XfQw2E/Z7jC0zzjvV4v
Wo3FOnwptnwX/U9y3HuXDmrovZWxfH9JpL7VoRcSOf8WwuE2W1PhimGuAczh5vr0
tyR27QKWEpOZcxMm/YXs3i82VJUvxDeuUjWGJYiO51+T0ZKPWK9HQ+q0sTqV84h/
C0bCs8CscMiZNcAZpjah1ACp0j4LrP0x+rJQqh+2rkLNs13dXQUjYCaU+4Rfy2Kc
wdd2FAtf9ALIGjt5xqTQaJz7DfkZ6UqYF4/OiY0zhHrk48FwqNPHi+uStceGy774
4wrUOGySpo5dAonzcvTiVL6oiU8cAShyq1I7+ksa7TnADgBXm3LxKEmlZ0Tg6LCn
ARNHicO45XXqWF95D2rR/BAp8/ESfL88WqKs4AcPPU9CgCgshCf8VOWg0Hodqlh7
BEy5r7S5snljw7nNmJh+mPjk5bkXSFH/NUY0BzZIVFAwgYn5LmE+cFGuAvsZ3Slf
8DGauon/3muoux4josr4Kf+/FqQ5ZV7sg14+lWva+b4wRp6ZUOlK0OzpAzNUoKOa
6Oh1PzH6gH7wBg0Hl5tp3KVhg/ZixrEt1Z1elDW0jweheiBGSOEHtfpftwXCU4EY
WHDok+lyJIqy77DUUZZp+lP9ABaL/VkHqvGQXhB3wWjm8FoYiN9SrRNChdy5E9Wg
Mzr2djZeicH5ID8QvlhsyTAbfVTrRwR+3MAU/8VZbvz1EbG8rj59RRB9Y9gPFmuK
NljNNx716FV54TcSPxhRDR4GySrHD5H9pgbjaz6g/2mVje84WQKL8MqsFpzLsvVW
0+7N3JJ8i+feLJVRKOS8+67QAC4K2MYlr1zene9xKk6CZ1EQO2Uvqqg0QSDMlbcU
Ykvezlix2xLQ2rea3tVh7I1NsPDPodMhobz1ZOTIp8BS+qBGL7K+CO2MQMoPCB+6
+jCrGZl7cH28daODPI3Q4R0wGDQCrwtEP89mpt16BLR7LFeP8kATALbQYt9hzjYj
bu6o2OjOMnoTsi+8u1EEfKmfgkGe9TFKjyWihtal/4e+MJZuTMKG+nNnD7nRtOTz
c0QM72hjEHntZDF84TLZenbSuQHqyOo/UD+k/3Kq2UfTmohy5yz8ik8Hbc/9zCeU
CzK52ym2IEvpqWgvUCvUQxX41Xx+Kfrs0FJ50H4BdLcoqYHv646qHW9KxR6zoSlo
0PoEs6lYW+dDWitsLvntbd5nmYdO/hTGTrGgUpxgXaWWBWM5RuEv+Y4A9Dd9vg0b
Cj7r3pl5C1LwmQy8OlQkkp+pNqpGu3lYYxmUgHyO1ehLKzY7zrEFnPYCruLZo7xG
EVy5np+v/yJCdThyXSb/vx0sbiXLJpojLRhTJSMilE9IXe8zYrPTmz3nUrNqLB1M
K7Mz1gumeKEslqGSkKLUV5mZ8zqxY8zEVI+rjf0/VxL98/cnEio4OVSHPTf73T9L
hVEk1ZNIuEFIYaqC5W6iKDhmKioAdzbFfEw9by+G3PqlWBD2W9byNN+ygdEH/qtV
ytEAt196PUJ/qFT5dm3n+5yumOwe1uYA7qj3Yw5vrPu7epMy9LnwqH9r3lL8ki77
+W8+PGLZ0NydU2zIX0tWWY2N2xVIvApW0SYE5PLkodWzBAywkeqDkv9Kpm8ebtPh
TRKafyt4EtFnBR9JD8Ka/hSeGe/sgbSFrLIoviwRn7Ala+HS6Qb6+z08JkGtRNYX
rI+TZN2dYb0jCNCyJpoP7f4q9dkuyFkHUoLoLgj8mzwBhlYz2W1aj2wimw2kEcj2
7wqIh0HfVAr7xFwzfd133Kegns+7IMV4duiTXJeYvDUrWi2KYb1KK/qxhTX6lUwb
vCl9XOjWrNbrZhkehycODzfjfF/GsqnYs3pO5zaJgzQr+ymRd5DVin3oB/77oZ+c
pLfBvYL93elm8Eee5azMRtroky4BaKgiFJwMLtC5aoT55cWa0W/vOKZFsvkLQ2ci
+hVUZLMNGMKhEcyTEA1B0UIaziqtOXZaMJJlw+BPWBfQqbhCE5Uw3EigGC20sZEc
rmfaOA/MWQbIUlgT4nU+LnVqUWhwqPNuN4zQ3UirMAyjZbTEgjmhyFpCKOA4dar+
7ostAzBscXqPIiR1G2jNne2Ynj1rYOmFNlVhO34zpZUIVOVST9bU/T4VA2h74942
tYGfMHXzS/d6NUTYnLh4uv95wjksXMWqKgKhIxA661RPUYUWJaRp9Vg7k2cc1+Wb
CWFoGfJFkEp2jJA7RmubzobSS2MrAyN4cEX9xUrnOqQeMcOnyyg1iGM6efqPWqqJ
uhUxV1ybrO54RsNsC0ZuxbPu8XzFfD/fFHjeP5/Zzd1luuJ4fB3Ne1oOoamqvTe7
a+zkh+o0IdqaMNWrC0siOXhLF5ZozDEJz0QfP3TMC1S+QY4fw647EeV5Gc8DBRq0
yAhPIgTH0lKPrp/4yV+FM9H9/hgI+xVZu55pfB90PwVaVYgWwBtuF3C9DE+3fGvN
iGrDkoOzWW5smY9UzKKWXSehMTxXIBQX24XGI+G+2Wqp+uyzFYT+jQzvQdJXsCu3
64+x+FHlA4cfNoHQKR52trTOv0Xt6X3svDF14rBkipvG4vsTdcZ5QH901jCRKmNc
cjAN2oSWVMkEzclocn7llGpSZlppwFT8+7/ZVrjxYD/xLpG9YAfqxG6cOOaw+dNz
O7DOKEm/OLLKnNctLapI/7Ycu1t1ch508zVlCNqcUncdvftD1bzR6X2UGgDWbOTd
9u9qQZHgHhUq4idyZidfICLrBPF+a7aKkLfg7nT4Jqmsl1GYaAOhxO4A/Q5oOLXg
EtjozcpG8YQzAbtPfaI5qRLkwqxxpzuMWkhLABz5JXcfj6uwvS9s61N9pnfBr41F
rISvnyVGVmZ2sDfLXiMH5v/yKn4lnYPkE+bJ/EvZOUoS1EXLzLrMaFNXbXWctE/M
fz4PETtkEg7338qKzetq1Tbgsnw8HAxJ2+F376XI9mR+bt44Nc4tSjj4KM4J3PwT
91okcwGvUns/QHqkLghMhRUtLYfPnibelwEniTvwJozBHGn1i0ky9KpsmsK3N8Rk
2jFGlTkRFfayqK84ZgiHNa7OwLiQ+BdfzSyEnjXQ4JFEZfysY5sfxZCDhv9BXkRw
bHtCH001MNSE7o3zW0pEYFTBjdvkJtFgpRwNO0HnTznxgtLP+/VCqlZU4Ko7SPyU
2s3+an4+t79Sg8jePxxMEYlgCWyTt5HAwkAR4scW7ur0kthgO5LjONnPTy81IDTo
EFWLih0GFppXFdt0tO28tyxl4Xe5N7jwN1laH3u62aT0WZkAAMG0pRztRkXXbBra
56wj8UpXP2kon8dvq5R3RRSwCoRnJ+D4FN2NMCYncxyB089D1RK+LsNKHWyE5AFZ
hKlk07T7q2w1LAzkA7h1dggmNIDCS/qNvVQXJuLULDNvphOsbwSxs9ICKVF6DZzd
gZSbUu7OVuW+MAe/YBiNTDYY0W8CUEUpz7MeUYCJmptFE9Ngssr6QREvDYUgU1pd
NPLxNY2EuB9IHKNIFPh0/lWermdhfcEN7Qb2onNTq0CkNFipAd6I2x10okbFJ0zh
pNW0CJxmqk08oro55WR/LHKLjnONFeWsOKCbgYD2LaqofiImI6CjY3ikB6q70IVv
44dVC5hrya28+hI+Hs9JOugSy7mqbSiowK9HdYodUiG5jlNYDAgahER7igYHDbHR
vHqCOMVWqTIAuCup54UHelrdmU7d6NUrgDsi7jT5fR3QegI9SM6Lx+upgIKiK+r7
4SVdHopFN3+yrRu1kidZAv868JmVcZQ72xFd1+r0RiHKTS5HA8ySKz0B5HwlZd81
0FvGlfbc4O7Lt5LpQQZEvdBoFBH/NoeI55Ky2fes5riPKBblaRUZnPIv2NHz3Twl
TSYcJrLG7zqmRQaevsnXHs4L/pwZPy5y6u+yHeD95n9ziW648lzMuSMoLeCdD+Z5
ShSeWFjDQzg9J1VtrfHwLKe5V6uJVEqnIwRb3l5EFqrqIO0VtQlMD7Idr4mpepkW
HLfz2hBIl9Fl1Fh/Piwvf3Xy9cTQZscOY9d5u49gFyNbc65qEu5i55SuRjPBzdcY
qii+32nC2/kguV/UbQYx9Zpq4Nt4gsEYS6iKrLqyG3Sk3yQYdkc11rfTkpe8bDdh
T7rC5vBt/OKMkgiH5OwP3Yo6/6CKNDAJ/2sqEITEUWRJjNOmbgXJ1DlZ3YiP4Hn7
aEpn+i33HKg2uCzdg/0LLLnuYXilqywxTghGEI/qtikPhnXkmxpqh3rx+B0dIOad
mQNYg/FHlJVdBzj9CSvRN5wc4EDFZ9ZYh/WQP6Ad3+Q8/xMlYUvG1LQ+4JbU347U
dQ7Ma8lq7ebiOmhckcnJ/wCERfXE/a3yeso0r2KXmT6jJw1nDmObmeNMcWuhun/r
BZV0frIm4vdIcERwAt1EjRyIuLIxpmt6OmoUpxqqMWZCLCZ1Ae4xpEZaquNw28qW
yeWEGfRiQqnXmueih/A8JNwQKZnGvG6BD7/3j9zNo1AzE8cmwAQW7DSvwx97SNFK
/M9lQmFhemEiXs91snDkkEeP/+bCZgJfrfLZUec5q0k9Yrr9M6gcvl1W00zL1C8h
8/jRQCf9XA+T0bgnmxcMbT27IWtSX9BvEFAofKrZXX+x1Mwt9tsWGep7h9AK0PE1
UarxWelG7APfi5whSKtPU1Qb9X6CvSrWiRHTY3XYDfexwqyssC6sfyak3VKf6W87
FHGCMSCt/OkkIY3mNP1wHMUOUzF4BtejwbkCo397SCLVJX9WrhF3wDxjlPH4JPNt
Pt2+6QJ6VYQfbiF53K+ijMT+Qzc6wtBllBI9vDErdQCSD7NWl6RxQC65NA51qUwG
9nyP1qBhLRdYtJDv+IT1JXiTs2odxoy+ykzCDjw++dO3dcx3GzAz7cwbDYy53TTg
rGkKr8zzxmp749TCAprHFHXYPtqaeOz/n+IWJIcTug3jNOicwAS/E5uazOAb7HDb
TxdIJC2c0TmoPqgEpryceXxNAN4aQi8V3V5ylAO10gpsDTY3GArCHpVEnxBoR57x
g+ZyQbfFDv4A5pxPRAB9jJSw54iF+QTHxBfpNSWn2ARfI6yWVjDzMs8dtSn61EWT
sMxh1PdDy8+MleUFemdku2aXsbhslfX+ODNX5x0DgEoA1eDTUH9K9HVTL2tZff89
dwaQErplYy6qIWUQ/18OnPeuw9w4WJ7PMG5meo4PyWYSj+alPJz3UMysz8sG30Of
zY/zYF+ennvsYfeEOriF0EUVylCYkM0XLxH2Cg2tSb8FZeDOkPRtxQaVJe7mFVIL
pzkVx5nbTuj3NGIV8qlcneXIw27kNqSOgG7STWqXg0vcJk4T7aBKQjhRrDzyS0FX
EVJvB+taQM1LDSorMaQKIgtyC3ErMavBQcTfFKBtaIMsJv1ACP6uV+4CbKCDdlmu
xMGBOPBoautsH6uqaO0S5LhEL1Nj9+wwu/E8+gXF+5ncFddpYyQGLajtaTqw+GY/
p6/fKUsxAnilmsrH44Ib8qUB+KaPeZ0AdgKpJu1U2rh7d/d6eo0gEKXTytkxorZw
o7fwuF+GLqSc7424nw05AQ/UrNnH7fluVZBhKwB/v+m51ET+7ThJXskz11ZZ6DNa
ei7Zff+fgyZba7BZDH75oRAdT6Qku0Fz2uL0awzpy1gpOQc2bLK2T/8SlGsIS5Tr
GoByrdbqY0rTJUB4qOgcqYNZMmE6qZMBlTOFb2zhgQCav1SG1fQ+i04jQGwrk9pI
cDbgvvYhAc2E+UZDDwiRyIyccgP/1TiEDp7feqfZK7S2PK5rnDjpd5Gf6PedHMPG
elCuWoi+dCarMaHHUIdGgEvRArzgeCMCa/2uAruF2Ln7XIo84r4qXbeSvp3IPspW
MgTcLsw+/tdmcdNzuU3AM9mVJG8Xq2XHy/WhOk0uV98k/KKAprHGSjLEoqB764zL
TV0VllNmpMGcJIOpMrxBga1D37jV1aaSVIwFVPa2V3Q7S5IiLawVjKnfXdLfKYn/
nNx0l8usBlpOVWc+flCSHUFbaaJO8zWv2EmetWjJg1coT0uSVPO9N40LifV41BnL
XEvn5wL2l2CLnnyjQEEdlGzkDcAybBw/z7Iop0n0lzunFPI0MRYhV6ayml7cGWds
FSrwt8WKI6iLZOVfcM+X+JWvRtyHlBi/C8aBd//BCBJjQnS+qN4e5/tUwXzH7kkI
zGWw5balAqXeIqDV0YMSSrLnUoL9hrM8lp5VGxKR4I6cL3dwtYhulITnwAZdzvUg
/bfSXPFYXmXIF5Z0DT0A0M0bTaWo0VXl1WiccMAvmAQ3hNy9oe1JXKMKyjnHBnYG
4AM+6JUI5j7lhFfTOHcwmJ20ll9TRqmb3JuuxSQ9pM1UJaS+ZWafkY+KwUhHW7kV
ORA3jZmDteRm2t6EKZsMsTDhBrymTu3N6pe8mRaCjJDSQysEHm+Mk++WixbnPGXq
mNH5Hh0ELiTLpqbsqPiBc/75ZOnHHlQBTzZ1bfOkjfzlcsM7sJTuiLqNekH6f6i0
AnydSet34Z6skO8f8t7VD+2aWtnxAGo/HwV0KCGnv0dTbmMqdYnveodibOgqn8iP
OXUJOsAQLq7zSKMjmSSJUWXMDXmJYE1feA3i6LQXfWShUnzhUDk+SDGsOoob3p42
dUKHDfSz37OHqORshIdQpvooJYwd1tOJTqjUwy/tk34QSrNo6k6DidprUqpOzaQ6
CA7oyZUjDyZy/dJiLRXrqFQNdGUlDku3bEiaTqP+xj29o0T1gLWeLfvIS8C6IzB5
77q5cyvw87Wbgx1313DePlRIlGPM/6FMzAu7dPPj+m7wOdwhSa82SIuTuwJLHyKo
ulpzZ/b4NRiYiPvu/VVzWjFEOsAg/FOmP8J0CDb6RP9ZqC3na1c1SfuRcPKookSH
l2CYS98ba8WnBu4HHoVBVpMr7NNv8Yuqrv4U/+O9Shf2vLDP+ZiB/sgYFglOlvlQ
ImdN4Eyudo5II+XS/IHXLXCmpNu3BV+IBQNde0hyM5N6WX9ZgR+2fte3Ks5REp65
tqwc2++IVV2h4+JpYr/D/YOp35jRul9GK2JEUC6+ik938Kg08cVbLeaN3+Qu7B58
EUwLFRpOAglHSxOozu/XIJgzUS3EORE64/hwhoJJXrKgybs5izkgsJelcUz0rQM2
m520iPngDzY+ZKxvRYLOeoSea/Fsi4Z3y+fJQbafX6v8z+0QMl2Fdfh3ZlrNZ1/C
Vdu1Id99e/Jso4RC/6AsTCjjENL/BtXPbeOsX5w74QyFtQKpnLTbmFxg5SnAnZ7Z
MtR6j4OmX9VmGg3Lb7q1LXlCfrpXmiV/C3YS3ioEt5Rz+COjuKwjlrIt3imBoKy3
M9FVpJg32xTUnGWaqWIgjBKLlUF5VwXhPig1SkSn53zkdDKr7O3zaljt0WFMUe3K
r7Mnn+dvi2kr2Pvby89CgX1kFKRMEA0l3vvYdzQhl2duhDsk/MMcuV1cMBTf5bli
+U4Z+S7Uwglm8yhjZTt513nH5o4Wl2XjVrbJK2+f95piAvYovwIHSMUupXtfgeEw
fmShlNEt8wE4M569ar0QIboXkasCJDfDlqmTJ30MEduxGQguhHVOTAbU3Qq4/T49
gU/0sWd/kUSIvluZnjMy/JpnuYA8IELGFjz74WFzsNZc79Gg9XR+lRdthgSn/231
/q+bNh0Tm00RtcDSZ/ugDkdtxOvqx1PmvTc2yNs1tRrRofhmZX1WVzN6iJ3pu2k1
NkXvxH1QrNoJmEGVgpJBonM8n+F7yr8fIvORiytWwDSM+xvEBgTU/39gVizeyIR1
d0GzrNbh7Iny0P8kzSQVqOnMSSfuIMrElyGZsQW12bmbSITqg9kpho0NXYoJau63
0iD8D+Bvi4hrprvoH0C6csSH283vGDIqOdbIULIRgTVFUmFtrnbq0s7Y6gd/Gwsj
4XQhNYaR475cTDt3k3ReAu9J5twKXedwjrGOf+ja1F7suRhbgSsYNCOFJat4JHMF
2XAS/4qF4fyf8jPMLGl/B1vpXHE1QDbm4VEy6NQE5KrA1NtoVjJtLvy9X0wVuyax
CP2X0NzF6VzS99GtEf+VAFQ+YJIfWAv/RUCIlU6PIH9MacnstVwUz+fvG4jd/gMW
BTy0JNE40oKMgwOXMTu3dMmysCb2uxWR37Tq3jvWCHHSCRPEHe2cH+AwIgZ9mwxa
hdigEpMnPAJQ4C4UWQThkYI0WyS5RoiGKLABsRdy0ulyX1NEDANjasxs4Y5bJ/Ll
xoFd0EJuJ7Rik7Dak/CAedzR4S7oFbsvvN3FXP3NwM6EqUThd4NSy/SN/FfvYQ7k
kC6tcYy3eEyoKL4q6MOJDnKiVHqqMgKgilm3Zhu43Whx7Jf59DGNeLwH91Ejimof
n3E0DZBlbClVo1PMecBgXVcZMs9CAhOGPDRkS/GmDHubtY2hbpKZlL0sL/GU4bRj
tLm/56WGyPAsxq6f22n3J+e83UTy37ZmiFnhaXUP9M6sP5yKPM3AzeK19PyEYxfy
PdZZr+FJamM6IRSw4z42zYK4VO7gKySxXZeBONt2QY7Lb2nTYY2+R/+0f4k4mOaC
hdhpNoOK8aKlszwlyRblfAx1xbAQYwY8YjQWNW3fHfgEX2iJHOGoUtQSb9Ur4aK1
ZxcyEhQ+sTQZV7NZB0FEp/o095FU3DGdG+IUtdL4kWRaK7dxmzenQ4B9jhg+r1Rs
M4C+G6iFVZunruzA027HMJxQFgQV7H0AJ8vhwgD29ht3YYPfrGjJzRja+ZPaiBwV
edzTxrPCBF93lxCh1sh5JKCYrnD758H6X/r4wxJ0gqjjjkn9YYbgRlhYshm2w6Cy
DmJHxfi8tZBZwPZC1WsMihJ5tV9rXnYb/2h9jJJVxe1LChWors7wOgZxQZsXArFh
aGtE0DOUQqtV/GNifJVNypZioBZEWrfN1fLXur3xbB723ccfEPQhGx/z3hqT2p/Q
UL4KXdhocUz68O55O5e2dR+6E2gq5VPhv36qHL7U/GGOKcf5rzj/Vm07C4DErkI4
lYUTo8LvA3/6l+gYrn4yOfy93F5Yy0SPnSwtrh4hXXklNmJ3D6NltUgYu8/rDha6
ewWJrI8zPxK/iwOaZRELIaiMse8ha9IHIc0mXM9H7nwD71FRLXgw3Ym4VQOzZM5z
OMJTNrjUsQOLw0zmtVsfGLBW3dt+ZWeBMSoZt/keATtBDVPD5WYUGEM6YyamzeGH
eHHQsAlpy1WmBr0myfemtK7/EzXngSZuSw158BY1gVjpnwvrMOpdnZP83RtYKbyb
/6D6YLILiiUetWups5neo9Ob99XPaTJd/VYy3Jz+9eyvkRP4/891spUej6koV8jR
hOwQsnzAAN1OfhfqjWTp5aupbF5zr7tjD5NxM/LLOnvYQ12x5qjJUxxKVtomIBSi
U/ADQOg+MOhD1X2bb0UlTTHw+ZVgYNqk5Zbaar3ADYsWedjNVtzviUwfK6B1LJbw
e8Oa6P6GWNNIZFeKuN3c+7fu9gSNGnrFma9215GJ+3j0u7/nK665ZIyX0MzmqUP7
0S00LfAT4SplGN4T1tX7KEm1CvE8FzikcylontBooGAMipdOCVZikRN24hqMsBj6
+b/hSuaLhAszsgccwQAugL+C/PJMm/pfS7wG1xHwNAAOt1HJNK9d4fnrUgo4RAOp
O6pGQbsi/H6b9/04W4pjbqQwz2bmdCQe+5O8ctQ5ASMYizmAMji/drHcZpXM110R
naBjFDlcQ1mZOXDAI3HBvwA1uCK1oorJXSY172/OoLki/cFVdgtE3xxemTsApqO7
B58FYykjCjwSKf3M3/LSK/0ta+9VJciogQzA2+vJBrnwurVrcY6JBuwcm6Gg6RCr
Zh5fZB+fTLfNQiaqZXFbVwLrd7D7BT/GoJiyiVutuwSWr3Maau8mSc8lrpQIHnjJ
IhC99rdP3OSDrRJqJ+ZEpMVTdkUsNRjpSXSpYcYpwr9wzUL8vmyPn/g3RM4r00de
QLve4FrUfVJLTIlzifQUYSWwdiZSfTwnK3GCqCYJUNon6qj7I9osbO0Tb0KmhUf3
VhUqW+P++nOYIOKNsfwV3EPiuP3DqTngP/xNrB8bsLt6UKdkBb9NnDkaGQiKTbO1
uSuxsO1Cdw86IOfIRWweamyfWamQF/1by4vcREe5dG8r03/iIpMJw2wnZ0VC7Zcy
CDNdfitVVY0/rCclJE6Ulrh0oSP4e0wds1v7qDc4T+ujmgSmshDkXFE1Slnhmp32
39mheJYKJBCFE8qN4YDazIZZhQLw+GjdZcO8jHhcU2wetcLE1QjKuZ+m1+AWJV9o
f+mec0ANEyT1g1YvVCAblEM1moPV2fHNS2+2ZF4UNlvuoGoZTc/pPGr4OnFr70Cq
38MUe8gTLEp+Ebi0MZBS55ATH3p18+JbJm7P9+CbZerB0eablbQR2HlfXrD4fpcn
FBythNiMFsF6udmikAAKioCoJ7Xa63s2jSFSbs8R8QdV9fxYekmC93WKWQO2fkkp
Nl4Bx0fAMILX8RWg7DFAFlw/YO0SrD/c1gJCa34n9jTyFa1mQKuqFgHotVgl7nsa
z5+KI6XJlXejMELbgdaXyuc9H6X22/2o1NpIBN2W9JJ/FTsh6DQ8sDI+75J4mZq3
oxTkjQuGOo9bzt9zXjrap+2I9S2cc4+tgS4IE7Sj6lkJqlKqdI6tEHuP4OcAfJvU
d5t6iEbssSRMPFb5IzVRiHD+noxyy2NJA2kxKH4ECvAk5LwHfx/gQSVlL4Jy6B9a
M6gOu6CIQaPqErYLYaNlSKcHEZ3xBolBtymBYkNArqokny5sZsGTkM1nVBQyzkCM
rQz6caZR6ZqEg/Ae/Ypqdb07O/48ZW8cyrZdvM+4suwDmd1kAsaGJ10xsazUNtsU
20iZyMAcvZ01BlUsxB9XZSllpUusdQh1O7OZz4qEDz/Dgd0RsLqZPukU/PLx6zK5
HS1hCQWiK/DZGpCZ6t0bjmj+4bjKP9pyrSBAG/k4dXykNM6m5PvsMI1x8vGOdJrC
wa7GD0vjgM9nm0enVXZqLNMe3KzcVhQ2ZVg8v3X/glapicvBqzhpfTO63a4LXWy4
ve8wZL++eIAlHDh+aZBM4oxWAh5Yt1u4mie6ejbHH0IUTgM53u6UdQCYW/jAk/8a
cMQZuWYhqf08GTUfJ5aC5EwYJoiI5t9hk5L2xzpxmSFhZHpq6jfDmhbC28tA29I1
BJ3D0cUTUpSALULX6fg6xQd3bc0EXcD94OJGMe6frBrSLHPPN/DsScqs3TyL+WZn
g7oPPeN+vOJRWNfFn4cu+vKeNClLGCr3P6qbQUOwotg0dGIg1cWpO0tvzoZUwIsM
tk52QgjApRAy4DyPA+1wCIWlJBWjxNnNNrbEGIlgFyEp23e6fg+ZSX7UJR5GE75O
ZkKwlwnwLuPkusd29nOhOzPZJT4iUSPwF74YSi4CAkh6vQHiJw2UBjNF21DCT4tr
a6kvD/yabzyCCuZJPQ3m+hY2FGpdQh+OUXRvmwQTauB0A36WZ+JxvCO9APs7TnxO
w0G4XFDTevTYpbYHM8TP+wRCTuElVHZ5GxTZxvRbibhnQOSYPay0CmdCSkwbBOSt
+x5+AOeB+p3BBIdUBvE6iAVKBubh9t8ONgCeQ39/Z1syZKdoxuULj9IX/QQ4qko1
41QBsvVjvFGy68R/ZJ9CCIoOiIfHMc57TDLHP/T70VXf0NDVs30QHRZpF2Va6LRR
uL1imo0hdDBEDx4jBa4SVw==
`pragma protect end_protected
