��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$��$�����Q�-E�zW�l5n$�0��4WO�G&z��|��T�<��r��Xz�q�*���*i�В-L_O�B��pL����V����d��Gc]%��u���c��D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&���~�`���sB��Zl�8&l���Q �h�/ޖ����1�L�-$|�v�����dϑ�"� u�ͣ��t��n�l_��?Y�E���>��;W��$�����H|�f(*�S��[9�
�c�^	��iǢ!m(5�����H�����@�LD��������w�����-B�B����>�"z)f�/��+!jtOk$ 4)ARBm�Bm5�|����sږ����ԢKdL�|��r��3����wN�J�ˡ�]W�/�)me�I���^��J
�j��̡J�uB�QFբ�ػ�$p~KA_�@jB=S����aPS���^s�7�2jS��4�o�h1���
U3�x?�-*ҷ��e会7�I>�*�{��|Ŋ�5~�N.��PU���lR )d_B��W�O�τ��x{��ݓ�i�z��W-ξ�E��IJ5��ʁ�M��,��.�m��h#��G��E��x\[`�� �����j�&c��BV��GSՅ�=�#օx�	�s��?1�|`#�8�y����kc�"i�/|Ӻ������|t|���7��aY����R~���8��:]���}�ze3}�uP��0ڱ��Tg<�<$��_��&�*M��k|�K�'��ґ���+��̩�/^��~�-�i��40��e����n�b�/PIo?��`o���R��{�7[E_�'� ���c�Gz�w�F���i��X0�Џ =	�m�e� �_��
H�L@��g�Q�iB���D�G֤�'�i��'9��n�K�)�3���'Yc������pO����Ey)��н瘶�᝟�/<w ��U�Ò�ܑ���Lԕ9@��b�	���_k��c�[؈���0�DhsD�ht��0[��_�]�x��BP�<�S���D�(����vy�P�i�?[�2P�A?`Y�o2���/��� �Q{Y�jd����D}6��A��0!�~ۜ�`�اְǲ�JXgP��T�X�\.��s�����L�=صe������'d�·Ư�)���_V��{9�U�� U���q�29�pꉅN_ZS����Z�y�Ҥ�: �`����@�M;M��Br$#�UT,�ޯj��G�톿{���a����>R{��!��!��2�{�Xk��W��S$J�t��$��sQ�1����W$:~�s��TƼl�0�e"]��'�&�����;���]�<�*���.�8��Ԧb������>��i���O<,g��F���򍓖�`h);Za�k��\즄k]1
��$	�R�Oq�5\7��s	�aU���DBk�4���f�+K����v����jb>�r޵C������NݑZ8[?d,x�� �����@�2������p��2�R5����إ�M�Ұ�M�q���n�����r���ާ2��Ѓ��	FB�����_�����]����]��7瘩�;ʋtm�4۠?��;w���@ԕ��&R�F����Im���9��M�VK�����'Y�����L���! ����>&�jugУ���V�i�N��4ظ�����M寧����/��Iv΁H<VTF���BAa?8�W���hm�Y,%��o#�S�b�G�4���2���$���
���S��i��"{HW����.!���%�t�-�������"2��,|��1��݃��[�8�؀� ���po����%������)#��)MZG$u���۔�ѭ���}݊���{=J�u��,�4X�&���t�g1D�b���U��Z7��|T�1l�-�/��n`3�9�M�%g���+��M4^L�����ȋ5��6�h���}l��$W?$��p�^��N	^(�0���.'�:𒨙�e�NwqM~B�c%Q����i�@I��e4�2�$Dv�2�*�����XC������Z^�7 ��2*2��A���#\xBk�CF�	tP��$^/��Gռ���o"2�;Z&	�lM���@"���rgVQ�c��gJ{�k�k/5-����ي{>�ؿ���l=5��t�#��
૸����a�l�CqP��0-B��cFl�@�2��A?��ha�CZ����v6Rꒁ��d�.:�'
���̮��W4�C���H\��t���?�N�`Ē��Ϋ��y��w?[���b�E0vy�*�sT<�3_!��$��'N���D�;�R������H����m����A�(�s��K���� ����ҏeU"9�?^�"�ܼ�N����ʅ���[G���B����G�o�Q��I� L�����p��}B<+�?�ņ����C8��$Łb��w�!!�MïGXY�/�32�*(l�٭�LR��8:{>%�*�Yb��sK�9���@َ�mSݞ5T0z�"y1&&
�o��f鋵Ful/P
u0�F�Б���[kh�R�_�a�ξ7V�Y�7�\���F�t��y�$��S��z#��)0�W���3�N6R!9���HޱV��~�r��詴Dz3���)���\I�?�.��]���<	�#J�h��Y����x�Ul��+��������ıM9WX�_�gH	�iG�+�Gb�#�hYEe-<�u�Xeew���Fh1(Y���G��@��>��!�����ݾ�ۑ�V�W��_�0g� ����\��?�'��D���V��-��C+��.u�<
@�����R�UI���
N����0�ut�n���$���WV��6�3�X�HqB�$���vA4��q�- B�\��?�w8!ɟC^�k�aGځ��E������p�	)������C#�CQ�3�9b�U��dÉ�n�� ���L¿�	6�i�3)�s_T��n�W�����Wc��v�+=Vt�vM%&�]�Eą���x�Z�����qsPV[W(��~:b �"�:�1�J*�&��A�I��tMY����m���+fz��4�˅������v��4�Z����t6?%��,��gR����V\�tf��b�@�[n�z��Ā���eD:�aږ�&[L�;]b��J����q�לFi��������0C&�iG�(P�o���O�^��E�}Eȉ�V��u�R����WD���+
�"PQ=BA�5�U�=�$IxV\"�}��ѣ��;:�Z���y���&��2n �|:����
�0W57t�=�FB�h�ɾ�a�?�A�ܲ�jp�c�T~�x� ��V �I���@٦��+^\ G)#�^�f��)A�V��q}
:�PlX����~*�	���h�2��⍚^�.m%�qY�%��UcJϜv�<PHfm���Pap��kgݥOcݕib�[R�q_�
����+��8>d��8g���B���2Ll��gm���]�2��-n�-�Kp�_�!<܊q���_��f��f��Qѯ0f�G��w>9������"�?Rֵ��X�JIP	Jm�f�>=��Q��G,�.3���L�������L�-U�`�:K����Mn�;�����4j���5+�� ����4\�7j'�6���V�R�ʬ�!�H�����r�@��H�^c��A\a!*"�����é��?�B�1邤�ݴ-V�J)���¨(-��E)ʸ���8z���9�|���� ��e�7�_)�Bٛof㝭�,�>�m7
��ة,~M`��Q��GU��ߔl�C3o��q�B]���XUb=�T����k�8&���R8��*��raC��Ь-'�b�C�,��\K��6r���$�S&s�?� B���d1���$��{	+z�/�At�0
ǧ�P�(-��Kh9E����'a�Y8�]1;�Nો45r�n<�)�eJ��	*3� [��1\�O���Qz�K��U!P�[m�3�RЏ}�� v��!��O�~/3:,l��qm��@=�hQ9��V��ɱ��v�����9�t��Jߚ#r(�}D�����SE���6Ѿ/xP�-K��S�
��}���!�%���yt��}�u�Ka<'L�܆�T#�B�Z8�U4&Ռ`{�s�9�m�xh2^��k�ql�h=.�m���Y�K�O��!�#ж%��l���d�/�+�Q�P]�#�D9[���@_v94��Ϗs�`���V���[�r�U�;�P������&X�)Z��*���V�M	I:��b���fxr�p�9eƺ�{`�/����.!��j�
���8�hh�����H�1���祷3WX-D��TH��q��Z��=*EIi��]���!���u[�1n"C� ���M@�z�vF�w�#�`�Q^�s=�| �[�2�R �0�1w��uDj��L?z��I���t�\R�O������ ����6�H�b���B[����:8��ْ<����X�;�bq��R�����1����2��v��F�<�ޅ��ϛs�{[��Y*/��00L=j�]ֆ�~�x7ׄ��*�v�6JUؙ����*?� Yjcm��U�Q��nV4IhY.7���DMB+U�t�����������b����]�a/U6؟�&��[0��ӣ�l��	���(�,B���GU7	��לH��boV�)��a�>"���d�*b[�p�H3>Ի�}�=��=����(��Usd�U��n�y�(�Q���*7T7����3rY��4�,i� {���W<2	�9|�if��3~�����D��UJ{�É��ܴn�>BǿL��)臚^;be %�k�j�_L�Vg�K��-��rp�_�Gup��դ���ݟHq����:���q��q
�ò�8Q��w�$⢓3�em�]x,Y���	6��#��zƤ���J���#�ߟw�A�H�U���N ���B���z�k�ߨ��	b���\�s����
.����K�[!�h���wʎH�śr�Q䋌n�H�f�]nX��g��W�3��y��qW�O�GQ��~� 9��)~�.Hk30e��k�\�Y��?����iu�ྺſo�>/�TY��sՁ�k��8�֨���ʭ����9>=�ڞt/�M�o8[3��ʦ�%1Pg� <�j�@��I�+A�8�����'lY�Oі�#�e�+�	��a��V��/<��E�PW1�J?��T֗�.}�R��MA�"]��q+H�?����E��H���C�l����jи	����Y9g'�ۂ٥c��D�ؚmURN�sTZ�9�7��P��P?�����@�7Q6hDR�fF�=�wh;� ��U�%����H�!�KqoM�hy)�C.U��^0�����%6*�e���� ��>�U�e0������u3n�zaz�*>��ψ��=�W���6`IJ
A�DW3g��H�)�Ճl��!��`U6Xc��uЉ鑚�%E�����8�������F�)"e ��GV֒�ܩ�����1��ʟ�K0Ncݼ 1�=����NKڮ:%߼u�wi�%�l�1<��=]fԷ���ϋR�iE�.�C,u{�cW��[��E�����}M���]{���a.bN��(���w��/�-}�,#��Y�D)E*w��?��c��^�&6��(���	�Ƃ��g���?�-M��.D�wa�d��`�{='��]��?�15�������|Wht�y��e����B(����Ş�m��E�밢��4���`�c[is��jNz{rc���E!gLm�8Pp�d���Rv��(�S����3[5{��;��s�������]rvw,jTz(���d��0n��X}�+��t�e��Ld Ty:��m������N$�_�n����ʚW�T�h���"�J���g�]?����|I)!��q��>$?����F�E�>�g������6�V	�-�}g�aD�,1���7l ��YT��MH�c���4w�͏� �䷁4�s7|9lR���]+�c���7��)r���{�Dʰ�7KG�WT�:WV�&9 �V/į�(��	/���v[<9hi_�V�S�rr@Ѷ��� �~	���xE�qz4R|F��&g�>;b��u�%��A����0��M�K�ݹ���v^�h`r�96b�Gҍ6���u���{��;�ğ3M�������j�j�ej㶼XH���&o�{���oXavڴ���Gd���`#ueoR�c�q�S&�L������-��&&wG�_W���(����%��B�l=(a�_�gsJ"4 ���N�V�NCV�ԄCn�ey}$SOIџ�z�OQ$������x
�'B��D1�|B$���ޭ�|���N��GR[��9�Mθj�U�a�+Ņ�ɛ�ac���ˋ���gmLU176�~ya�����Ͳ}(�/�Q�Lﱊ�@�C�zI��VO�:�7��k.o\�`?�э�z�;�S�
�[��@�a�?����ă)lpF��ވ&۱Њ~�+4��F�9�0� ��`��6u�\m[33E�9�z�9��9��$�D����Z����S}���*��e�u(�9�Ir�6n��P�a߮SP��l�'��xy�m�@�ƣ.�oi�+c� � ����3M�O�H,g�h��tϒ��o�d����Aq�[�q\&thA��
6BVfj��E���qUHD�A���I��O����2��e�H�Û�y�'�4>3��t�D��k��ʽ�e8�@��F���y�[%�����}$U:דd�3$�N��r��ީ����LO,>�=��^��Ce��*Y�?T�eM"���7�us��-�F��e���c�q�4�v�	��9��o�� w���7��sO."�9��~I���w诬w�E�}��=�;�&�Z<ة-�9���\�ɭ"����3xN���h&gڶ�#߻��V�Y�u6��ž�/[�g���|���E�pT!.�g��6�::�	@������h��"G���Փ;�[tڮ�b/����ŭ�d�����θZ��л�G�}C�@B���`I�~�Դ���^oWȡ&	�C�ɇ��I'8�=`��N֏�+��x�܃ȝ �i�p�ـE*��8��d'좨�D����nz���}ၕ)���ho�:�c!w4��L�q�zf�@>nn!��q��M^u��!�|+��a��w��=V���5R��ٟ������F�T�-'JK��������Is�g*�b��CG�c ��>g�tE�$M}x���M.!�[�6~���?��o�IQ�[���K�~�DF�-Ξa���\����g�w��T�Oۿ�4�T�k�cωq>O���yߝ���~�L���77f�e�ؾ��Wgm<ZJ��.�<G�X�R�}��#$p$L`4qy�r燅�T�!��Z�m6�`�{��+깱/|��f���+y�N5�����q�5���Њo�.^V�-,1�2���]��O��I�[�MQ���K��\߅)lv���Y�DF*u�̍��^C��?��n	�k�/h`�{����g��#�-Ga�1�� $ȷ5f���
o��ӫ� ���'����öw���+_�]H[�jP]"����m��@8�q@1�;�xş`�)c�o(�����z��j�$rz�o���;.�Z�ӹ����U�m?..��Ba�)�ѵ�Њ�C�~zX!
)�MW�	Hil�UhqP��-��f�dV��SD!���{�"[����p~��[:t�y:���;T�N�sD
`�vr+;�WY�d�j�+ԴQ-�Y����u��2�-r����ow@"�����i-l�x!mU Wa`"ơ�r6B���3_|�����$�xL�b���/�l�s�%E��x~x{�x1V�0w�R�k���)	���Ť��ސ.����VF��fZUk��K���g�k��F��h�:$�F߅��_��9G��M/8��d���m�o�˗�To�؏��O/g���8t\�<,���4�G��]d\�1�\�&��{�z/6��2d$/O3�[���\n%�������M��G�&���6a�<����0������+���X/�p�I4�}
E<��$)������U3+um�oU\�[�׊�H����7d�AblKKP��*��j�*���{rW����Bd-3��x/9���~��N3���:�M�U��7r�V��Qo��hC�t33�M��x�����sZ�"dI�k!������<(��;�fB�Z);U)�`'�3*!��k�KQJ,�sζ��*�.-�Ҵ� W�~��HG@��*=��'��x+��
�weET��N'��0�߅��@�=�@���O]���_�)�!A��Cg��ٹa�����T*N��^��f�nŲ��!�@1�����Ҋ$@Zo��[�Ҁ�Ғ7��8����-M.L�dw���"n����?F���,`��+�2���D^�i�H���Kҝrr���]ھK������x��É�vȒ��<���!,p����]6�1�;X���Eu�R:	аp��JbX샃e�2�X��r3E�1�N���^��/��{��һT|�1�!�Nx��Zs�Z���.�3+}�g�I9'�v;��P m�mY��8��1s�j>5������^�Ã5��9�%�	���Ar�h�g�z�R2;a	_��wI�������u�mB�����u��Ε�_/�oU��T⩺�ى��GG�0��fz���eԠ�|��*8�|�C� A�&4��d^j��t�꾆,^�`�v��C��{�W��?.8;Ӈ������.2�s���YO�;V��WfIv���5�雠�t�g9��ɥ]�\RZ�VL���Em�.>[�0�uP?��]NM����*ae��MБ ?��R��u��`�}�Vf�#��t�v��+�f�@D@�ܡ�'�to�5j��$�QP&����M;��o�!�@�N��-��|��̈[Mm�6�������:كgƧjտ^/�R�V��dB�����-�&H rOˬ6#sx��ӎ��v�7�Ό��nxV��G�7�����D)@�]	Bl����.��������3!�^��$M�j�r؟\�/a����ȋf�W����^n
�� ��=VP�!���&�B}��:P=\h|H�۳O�魯��
<{ۦd8�0~��W-��߱"d���B%�PQ��؉�3\�+>ز�?B9Īx��
N[I��n
 ^�sʤB\N"�(%�P}@}��M�=;�R�xs(�
1�3y�Mu���$������#P`
k��3`��ߎi�pK>Pkk��&yc�O��h��H�e�+5Gr?��/���u��<��[{I���'��*y�)����/Ut�R��Ⱥ����`�Kq
�wը-�p9�h*f.k�<��2�4*W~��.?��y�S����(�u��_,��U�l#Z		o<�Y{>v^Z(�����k�w�g� ;���C��qD1(���m/#J\��mL�&�v��	�V��W��u%�35'NhB�u'����R��CXJ��D�,�Vh:ұ��|q7m�CI�L�;�_�7�{��֮�n�v��փݚ�P2@OI{8��oV�t�&�)c�M�$�o�V.�&5��>eJ�n�|���7$�; ������5�Os������;=�;�Mtւ���qd�T��p>)�Hd7)���X4S���Q�7±ف�*ŝ�[���u#9Qor����;"t��3��ڄj�V8�a�H����'O�E�whA]n���*$�Z���<l��d>�	����Sl�S�^'��K�\���v��;�4��+�.� Z�R��̈�����۴X]��B�Zt�a���]2�7�=��{�lX
a��H��<QҀ�r��}���=��YN�L�k *�����P
g��Tg����+G��zSk�c�~` aǍ�d!9�bP6�:ٷZ0�{����իo��ʕ�7�]Z��$Kؓ�������H���~�%u���C'hVza��5�Έ<j�	���"����ݦ�_C[)�m��w���qd0��q)�>�Y�f��CW|� Z�l9䇪[^�����Z��[sf@G k�Z��Tŗ���Ӊ$ʴq��x�A-�@j�ek9�d[b.0�X��F,�d�B`�Q�c(eu���ܒ`�1���@)JB| �z��R��L�P>�"#����`�O|~����Û���@�����O!�6����FΔ�G)�uR�	�?-�>�|���v�ٗ��'����CL���:���LP*�B�����Wt�"?���Xtp}qQ��q�������p|ԻUOoY��ur�,��Gyʫ�!�vp�alo^V��nTL��ۮ��Z7�-��d� �Ȃ�A��=��=�/{���w�e��E#=��[Y2�+^��e2$Y��P��}�q�5i��(�~�[{�0�Q�xM{�O�a{��\�2K�^F�v_�q����,��|'�N?bp������;gW��$PDve���xFࣧ��jL�er_���J/����=:�p�
��� �Y�a��ʻ�#z6l����_�n�LV1m�e���R7Z�T(v�����4�8$�ΰ��Ý�Z,T��Ps�]%��0+����ϛ�w���-wMM��yHf��e�ì��o��\�; ��%f%�D�pG�0Q�t���'Yݒ{�B�����7J�}�W�m N�W���<4�)67�몖���Eҧ�r�V'<E�:d�R��x�wYШ���b/�nRБ��i��8ԁ!�l�G�s��Ԓ��遨��ҝ�����������+���.�Y��oH����"�S�x��kv=�R�NB6�����+�4�erܨ���JFPY�~�u�AO�|�?��!  ��Q�o;"�h�>�W��""U'�L������&�����ww���G��4R�A(��*�k�e� ������Ӄ��b[LD���Q��C̀�S޿)��b�R���Ռ�_�(�f}�O�� z�����66� �%_�7�@y��Kl����F�y�diy��D7��]��ȯ��PӼ+��v1�΃�;��{�~ ��)��-[I �K� ��c��]\!�2(fO29���Tg���%��6L|���A��\�P�I�}��7��3�v�X�y�K8ϔ�����cP8��.F�<]� ~zٰ�R�$Q�N�|��*��о9*9�֔�z��K㳗?�ғy��U7�嗲�dL��ڀ./'��dk̩�+ItZR�3�l�E��75z+���SV7<�~]��J*T��/w�~��H�-E��fNQ�w��o��QI���"� �
(���>4�j�^�����PJ�O<ˬ�_-�"���:���1�3)��`K�~��'���3�4�(�